----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 02/16/2022 05:11:46 PM
-- Design Name: 
-- Module Name: mpg - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity mpg is
    Port ( en : out STD_LOGIC;
           input : in STD_LOGIC;
           clock : in STD_LOGIC);
end mpg;

architecture Behavioral of mpg is

signal count_int : std_logic_vector(15 downto 0) :=x"0000";
signal Q1 : std_logic :='0';
signal Q2 : std_logic :='0';
signal Q3 : std_logic :='0';

begin

en <= Q2 AND (NOT Q3);

process(clock)
begin
    if clock'event and clock='1' then
        count_int <= count_int + 1;
    end if;
end process;

process(clock)
begin
    if clock'event and clock='1' then
        if count_int = "1111111111111111" then
            Q1 <= input;
        end if;
    end if;
end process;

process(clock)
begin
    if clock'event and clock='1' then
        Q2 <= Q1;
        Q3 <= Q2;
    end if;
end process;

end Behavioral;
